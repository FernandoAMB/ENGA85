// medidor_desempenho.v

// Generated using ACDS version 17.1 590

`timescale 1 ps / 1 ps
module medidor_desempenho (
		input  wire        clk_clk,             //        clk.clk
		output wire [31:0] clockcount_readdata, // clockcount.readdata
		input  wire        reset_reset_n,       //      reset.reset_n
		output wire [31:0] sum_readdata         //        sum.readdata
	);

	wire  [31:0] nios2_qsys_0_data_master_readdata;                                  // mm_interconnect_0:nios2_qsys_0_data_master_readdata -> nios2_qsys_0:d_readdata
	wire         nios2_qsys_0_data_master_waitrequest;                               // mm_interconnect_0:nios2_qsys_0_data_master_waitrequest -> nios2_qsys_0:d_waitrequest
	wire         nios2_qsys_0_data_master_debugaccess;                               // nios2_qsys_0:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_qsys_0_data_master_debugaccess
	wire  [16:0] nios2_qsys_0_data_master_address;                                   // nios2_qsys_0:d_address -> mm_interconnect_0:nios2_qsys_0_data_master_address
	wire   [3:0] nios2_qsys_0_data_master_byteenable;                                // nios2_qsys_0:d_byteenable -> mm_interconnect_0:nios2_qsys_0_data_master_byteenable
	wire         nios2_qsys_0_data_master_read;                                      // nios2_qsys_0:d_read -> mm_interconnect_0:nios2_qsys_0_data_master_read
	wire         nios2_qsys_0_data_master_write;                                     // nios2_qsys_0:d_write -> mm_interconnect_0:nios2_qsys_0_data_master_write
	wire  [31:0] nios2_qsys_0_data_master_writedata;                                 // nios2_qsys_0:d_writedata -> mm_interconnect_0:nios2_qsys_0_data_master_writedata
	wire  [31:0] nios2_qsys_0_instruction_master_readdata;                           // mm_interconnect_0:nios2_qsys_0_instruction_master_readdata -> nios2_qsys_0:i_readdata
	wire         nios2_qsys_0_instruction_master_waitrequest;                        // mm_interconnect_0:nios2_qsys_0_instruction_master_waitrequest -> nios2_qsys_0:i_waitrequest
	wire  [16:0] nios2_qsys_0_instruction_master_address;                            // nios2_qsys_0:i_address -> mm_interconnect_0:nios2_qsys_0_instruction_master_address
	wire         nios2_qsys_0_instruction_master_read;                               // nios2_qsys_0:i_read -> mm_interconnect_0:nios2_qsys_0_instruction_master_read
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect;         // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata;           // jtag_uart_0:av_readdata -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest;        // jtag_uart_0:av_waitrequest -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address;            // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read;               // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_read -> jtag_uart_0:av_read_n
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write;              // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_write -> jtag_uart_0:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata;          // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	wire  [31:0] mm_interconnect_0_acumulador_0_avalon_slave_0_readdata;             // Acumulador_0:readdata -> mm_interconnect_0:Acumulador_0_avalon_slave_0_readdata
	wire         mm_interconnect_0_acumulador_0_avalon_slave_0_read;                 // mm_interconnect_0:Acumulador_0_avalon_slave_0_read -> Acumulador_0:read
	wire         mm_interconnect_0_acumulador_0_avalon_slave_0_write;                // mm_interconnect_0:Acumulador_0_avalon_slave_0_write -> Acumulador_0:write
	wire  [31:0] mm_interconnect_0_acumulador_0_avalon_slave_0_writedata;            // mm_interconnect_0:Acumulador_0_avalon_slave_0_writedata -> Acumulador_0:writedata
	wire  [31:0] mm_interconnect_0_medidor_de_desempenho_0_avalon_slave_0_readdata;  // Medidor_de_Desempenho_0:readdata -> mm_interconnect_0:Medidor_de_Desempenho_0_avalon_slave_0_readdata
	wire         mm_interconnect_0_medidor_de_desempenho_0_avalon_slave_0_read;      // mm_interconnect_0:Medidor_de_Desempenho_0_avalon_slave_0_read -> Medidor_de_Desempenho_0:read
	wire         mm_interconnect_0_medidor_de_desempenho_0_avalon_slave_0_write;     // mm_interconnect_0:Medidor_de_Desempenho_0_avalon_slave_0_write -> Medidor_de_Desempenho_0:write
	wire  [31:0] mm_interconnect_0_medidor_de_desempenho_0_avalon_slave_0_writedata; // mm_interconnect_0:Medidor_de_Desempenho_0_avalon_slave_0_writedata -> Medidor_de_Desempenho_0:writedata
	wire  [31:0] mm_interconnect_0_nios2_qsys_0_debug_mem_slave_readdata;            // nios2_qsys_0:debug_mem_slave_readdata -> mm_interconnect_0:nios2_qsys_0_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios2_qsys_0_debug_mem_slave_waitrequest;         // nios2_qsys_0:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_qsys_0_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios2_qsys_0_debug_mem_slave_debugaccess;         // mm_interconnect_0:nios2_qsys_0_debug_mem_slave_debugaccess -> nios2_qsys_0:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios2_qsys_0_debug_mem_slave_address;             // mm_interconnect_0:nios2_qsys_0_debug_mem_slave_address -> nios2_qsys_0:debug_mem_slave_address
	wire         mm_interconnect_0_nios2_qsys_0_debug_mem_slave_read;                // mm_interconnect_0:nios2_qsys_0_debug_mem_slave_read -> nios2_qsys_0:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios2_qsys_0_debug_mem_slave_byteenable;          // mm_interconnect_0:nios2_qsys_0_debug_mem_slave_byteenable -> nios2_qsys_0:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios2_qsys_0_debug_mem_slave_write;               // mm_interconnect_0:nios2_qsys_0_debug_mem_slave_write -> nios2_qsys_0:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios2_qsys_0_debug_mem_slave_writedata;           // mm_interconnect_0:nios2_qsys_0_debug_mem_slave_writedata -> nios2_qsys_0:debug_mem_slave_writedata
	wire         mm_interconnect_0_data_memory_s1_chipselect;                        // mm_interconnect_0:data_memory_s1_chipselect -> data_memory:chipselect
	wire  [31:0] mm_interconnect_0_data_memory_s1_readdata;                          // data_memory:readdata -> mm_interconnect_0:data_memory_s1_readdata
	wire  [10:0] mm_interconnect_0_data_memory_s1_address;                           // mm_interconnect_0:data_memory_s1_address -> data_memory:address
	wire   [3:0] mm_interconnect_0_data_memory_s1_byteenable;                        // mm_interconnect_0:data_memory_s1_byteenable -> data_memory:byteenable
	wire         mm_interconnect_0_data_memory_s1_write;                             // mm_interconnect_0:data_memory_s1_write -> data_memory:write
	wire  [31:0] mm_interconnect_0_data_memory_s1_writedata;                         // mm_interconnect_0:data_memory_s1_writedata -> data_memory:writedata
	wire         mm_interconnect_0_data_memory_s1_clken;                             // mm_interconnect_0:data_memory_s1_clken -> data_memory:clken
	wire         mm_interconnect_0_program_memory_s1_chipselect;                     // mm_interconnect_0:program_memory_s1_chipselect -> program_memory:chipselect
	wire  [31:0] mm_interconnect_0_program_memory_s1_readdata;                       // program_memory:readdata -> mm_interconnect_0:program_memory_s1_readdata
	wire  [12:0] mm_interconnect_0_program_memory_s1_address;                        // mm_interconnect_0:program_memory_s1_address -> program_memory:address
	wire   [3:0] mm_interconnect_0_program_memory_s1_byteenable;                     // mm_interconnect_0:program_memory_s1_byteenable -> program_memory:byteenable
	wire         mm_interconnect_0_program_memory_s1_write;                          // mm_interconnect_0:program_memory_s1_write -> program_memory:write
	wire  [31:0] mm_interconnect_0_program_memory_s1_writedata;                      // mm_interconnect_0:program_memory_s1_writedata -> program_memory:writedata
	wire         mm_interconnect_0_program_memory_s1_clken;                          // mm_interconnect_0:program_memory_s1_clken -> program_memory:clken
	wire         irq_mapper_receiver0_irq;                                           // jtag_uart_0:av_irq -> irq_mapper:receiver0_irq
	wire  [31:0] nios2_qsys_0_irq_irq;                                               // irq_mapper:sender_irq -> nios2_qsys_0:irq
	wire         rst_controller_reset_out_reset;                                     // rst_controller:reset_out -> [Acumulador_0:reset_n, mm_interconnect_0:Acumulador_0_reset_reset_bridge_in_reset_reset]
	wire         rst_controller_001_reset_out_reset;                                 // rst_controller_001:reset_out -> [Medidor_de_Desempenho_0:reset_n, data_memory:reset, irq_mapper:reset, jtag_uart_0:rst_n, mm_interconnect_0:nios2_qsys_0_reset_reset_bridge_in_reset_reset, nios2_qsys_0:reset_n, program_memory:reset, rst_translator:in_reset]
	wire         rst_controller_001_reset_out_reset_req;                             // rst_controller_001:reset_req -> [data_memory:reset_req, nios2_qsys_0:reset_req, program_memory:reset_req, rst_translator:reset_req_in]
	wire         nios2_qsys_0_debug_reset_request_reset;                             // nios2_qsys_0:debug_reset_request -> rst_controller_001:reset_in1

	Acumulador_Interface acumulador_0 (
		.reset_n    (~rst_controller_reset_out_reset),                         //          reset.reset_n
		.write      (mm_interconnect_0_acumulador_0_avalon_slave_0_write),     // avalon_slave_0.write
		.writedata  (mm_interconnect_0_acumulador_0_avalon_slave_0_writedata), //               .writedata
		.read       (mm_interconnect_0_acumulador_0_avalon_slave_0_read),      //               .read
		.readdata   (mm_interconnect_0_acumulador_0_avalon_slave_0_readdata),  //               .readdata
		.sum_export (sum_readdata),                                            //    conduit_end.readdata
		.clock      (clk_clk)                                                  //          clock.clk
	);

	clockCounter medidor_de_desempenho_0 (
		.reset_n      (~rst_controller_001_reset_out_reset),                                //          reset.reset_n
		.read         (mm_interconnect_0_medidor_de_desempenho_0_avalon_slave_0_read),      // avalon_slave_0.read
		.write        (mm_interconnect_0_medidor_de_desempenho_0_avalon_slave_0_write),     //               .write
		.writedata    (mm_interconnect_0_medidor_de_desempenho_0_avalon_slave_0_writedata), //               .writedata
		.readdata     (mm_interconnect_0_medidor_de_desempenho_0_avalon_slave_0_readdata),  //               .readdata
		.extern_count (clockcount_readdata),                                                //    conduit_end.readdata
		.clock        (clk_clk)                                                             //          clock.clk
	);

	medidor_desempenho_data_memory data_memory (
		.clk        (clk_clk),                                     //   clk1.clk
		.address    (mm_interconnect_0_data_memory_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_data_memory_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_data_memory_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_data_memory_s1_write),      //       .write
		.readdata   (mm_interconnect_0_data_memory_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_data_memory_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_data_memory_s1_byteenable), //       .byteenable
		.reset      (rst_controller_001_reset_out_reset),          // reset1.reset
		.reset_req  (rst_controller_001_reset_out_reset_req),      //       .reset_req
		.freeze     (1'b0)                                         // (terminated)
	);

	medidor_desempenho_jtag_uart_0 jtag_uart_0 (
		.clk            (clk_clk),                                                     //               clk.clk
		.rst_n          (~rst_controller_001_reset_out_reset),                         //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                     //               irq.irq
	);

	medidor_desempenho_nios2_qsys_0 nios2_qsys_0 (
		.clk                                 (clk_clk),                                                    //                       clk.clk
		.reset_n                             (~rst_controller_001_reset_out_reset),                        //                     reset.reset_n
		.reset_req                           (rst_controller_001_reset_out_reset_req),                     //                          .reset_req
		.d_address                           (nios2_qsys_0_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios2_qsys_0_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios2_qsys_0_data_master_read),                              //                          .read
		.d_readdata                          (nios2_qsys_0_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios2_qsys_0_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios2_qsys_0_data_master_write),                             //                          .write
		.d_writedata                         (nios2_qsys_0_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (nios2_qsys_0_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios2_qsys_0_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios2_qsys_0_instruction_master_read),                       //                          .read
		.i_readdata                          (nios2_qsys_0_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios2_qsys_0_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (nios2_qsys_0_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (nios2_qsys_0_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios2_qsys_0_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios2_qsys_0_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios2_qsys_0_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios2_qsys_0_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios2_qsys_0_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios2_qsys_0_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios2_qsys_0_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios2_qsys_0_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                            // custom_instruction_master.readra
	);

	medidor_desempenho_program_memory program_memory (
		.clk        (clk_clk),                                        //   clk1.clk
		.address    (mm_interconnect_0_program_memory_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_program_memory_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_program_memory_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_program_memory_s1_write),      //       .write
		.readdata   (mm_interconnect_0_program_memory_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_program_memory_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_program_memory_s1_byteenable), //       .byteenable
		.reset      (rst_controller_001_reset_out_reset),             // reset1.reset
		.reset_req  (rst_controller_001_reset_out_reset_req),         //       .reset_req
		.freeze     (1'b0)                                            // (terminated)
	);

	medidor_desempenho_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                                    (clk_clk),                                                            //                                clk_0_clk.clk
		.Acumulador_0_reset_reset_bridge_in_reset_reset   (rst_controller_reset_out_reset),                                     // Acumulador_0_reset_reset_bridge_in_reset.reset
		.nios2_qsys_0_reset_reset_bridge_in_reset_reset   (rst_controller_001_reset_out_reset),                                 // nios2_qsys_0_reset_reset_bridge_in_reset.reset
		.nios2_qsys_0_data_master_address                 (nios2_qsys_0_data_master_address),                                   //                 nios2_qsys_0_data_master.address
		.nios2_qsys_0_data_master_waitrequest             (nios2_qsys_0_data_master_waitrequest),                               //                                         .waitrequest
		.nios2_qsys_0_data_master_byteenable              (nios2_qsys_0_data_master_byteenable),                                //                                         .byteenable
		.nios2_qsys_0_data_master_read                    (nios2_qsys_0_data_master_read),                                      //                                         .read
		.nios2_qsys_0_data_master_readdata                (nios2_qsys_0_data_master_readdata),                                  //                                         .readdata
		.nios2_qsys_0_data_master_write                   (nios2_qsys_0_data_master_write),                                     //                                         .write
		.nios2_qsys_0_data_master_writedata               (nios2_qsys_0_data_master_writedata),                                 //                                         .writedata
		.nios2_qsys_0_data_master_debugaccess             (nios2_qsys_0_data_master_debugaccess),                               //                                         .debugaccess
		.nios2_qsys_0_instruction_master_address          (nios2_qsys_0_instruction_master_address),                            //          nios2_qsys_0_instruction_master.address
		.nios2_qsys_0_instruction_master_waitrequest      (nios2_qsys_0_instruction_master_waitrequest),                        //                                         .waitrequest
		.nios2_qsys_0_instruction_master_read             (nios2_qsys_0_instruction_master_read),                               //                                         .read
		.nios2_qsys_0_instruction_master_readdata         (nios2_qsys_0_instruction_master_readdata),                           //                                         .readdata
		.Acumulador_0_avalon_slave_0_write                (mm_interconnect_0_acumulador_0_avalon_slave_0_write),                //              Acumulador_0_avalon_slave_0.write
		.Acumulador_0_avalon_slave_0_read                 (mm_interconnect_0_acumulador_0_avalon_slave_0_read),                 //                                         .read
		.Acumulador_0_avalon_slave_0_readdata             (mm_interconnect_0_acumulador_0_avalon_slave_0_readdata),             //                                         .readdata
		.Acumulador_0_avalon_slave_0_writedata            (mm_interconnect_0_acumulador_0_avalon_slave_0_writedata),            //                                         .writedata
		.data_memory_s1_address                           (mm_interconnect_0_data_memory_s1_address),                           //                           data_memory_s1.address
		.data_memory_s1_write                             (mm_interconnect_0_data_memory_s1_write),                             //                                         .write
		.data_memory_s1_readdata                          (mm_interconnect_0_data_memory_s1_readdata),                          //                                         .readdata
		.data_memory_s1_writedata                         (mm_interconnect_0_data_memory_s1_writedata),                         //                                         .writedata
		.data_memory_s1_byteenable                        (mm_interconnect_0_data_memory_s1_byteenable),                        //                                         .byteenable
		.data_memory_s1_chipselect                        (mm_interconnect_0_data_memory_s1_chipselect),                        //                                         .chipselect
		.data_memory_s1_clken                             (mm_interconnect_0_data_memory_s1_clken),                             //                                         .clken
		.jtag_uart_0_avalon_jtag_slave_address            (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),            //            jtag_uart_0_avalon_jtag_slave.address
		.jtag_uart_0_avalon_jtag_slave_write              (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),              //                                         .write
		.jtag_uart_0_avalon_jtag_slave_read               (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),               //                                         .read
		.jtag_uart_0_avalon_jtag_slave_readdata           (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),           //                                         .readdata
		.jtag_uart_0_avalon_jtag_slave_writedata          (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),          //                                         .writedata
		.jtag_uart_0_avalon_jtag_slave_waitrequest        (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest),        //                                         .waitrequest
		.jtag_uart_0_avalon_jtag_slave_chipselect         (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),         //                                         .chipselect
		.Medidor_de_Desempenho_0_avalon_slave_0_write     (mm_interconnect_0_medidor_de_desempenho_0_avalon_slave_0_write),     //   Medidor_de_Desempenho_0_avalon_slave_0.write
		.Medidor_de_Desempenho_0_avalon_slave_0_read      (mm_interconnect_0_medidor_de_desempenho_0_avalon_slave_0_read),      //                                         .read
		.Medidor_de_Desempenho_0_avalon_slave_0_readdata  (mm_interconnect_0_medidor_de_desempenho_0_avalon_slave_0_readdata),  //                                         .readdata
		.Medidor_de_Desempenho_0_avalon_slave_0_writedata (mm_interconnect_0_medidor_de_desempenho_0_avalon_slave_0_writedata), //                                         .writedata
		.nios2_qsys_0_debug_mem_slave_address             (mm_interconnect_0_nios2_qsys_0_debug_mem_slave_address),             //             nios2_qsys_0_debug_mem_slave.address
		.nios2_qsys_0_debug_mem_slave_write               (mm_interconnect_0_nios2_qsys_0_debug_mem_slave_write),               //                                         .write
		.nios2_qsys_0_debug_mem_slave_read                (mm_interconnect_0_nios2_qsys_0_debug_mem_slave_read),                //                                         .read
		.nios2_qsys_0_debug_mem_slave_readdata            (mm_interconnect_0_nios2_qsys_0_debug_mem_slave_readdata),            //                                         .readdata
		.nios2_qsys_0_debug_mem_slave_writedata           (mm_interconnect_0_nios2_qsys_0_debug_mem_slave_writedata),           //                                         .writedata
		.nios2_qsys_0_debug_mem_slave_byteenable          (mm_interconnect_0_nios2_qsys_0_debug_mem_slave_byteenable),          //                                         .byteenable
		.nios2_qsys_0_debug_mem_slave_waitrequest         (mm_interconnect_0_nios2_qsys_0_debug_mem_slave_waitrequest),         //                                         .waitrequest
		.nios2_qsys_0_debug_mem_slave_debugaccess         (mm_interconnect_0_nios2_qsys_0_debug_mem_slave_debugaccess),         //                                         .debugaccess
		.program_memory_s1_address                        (mm_interconnect_0_program_memory_s1_address),                        //                        program_memory_s1.address
		.program_memory_s1_write                          (mm_interconnect_0_program_memory_s1_write),                          //                                         .write
		.program_memory_s1_readdata                       (mm_interconnect_0_program_memory_s1_readdata),                       //                                         .readdata
		.program_memory_s1_writedata                      (mm_interconnect_0_program_memory_s1_writedata),                      //                                         .writedata
		.program_memory_s1_byteenable                     (mm_interconnect_0_program_memory_s1_byteenable),                     //                                         .byteenable
		.program_memory_s1_chipselect                     (mm_interconnect_0_program_memory_s1_chipselect),                     //                                         .chipselect
		.program_memory_s1_clken                          (mm_interconnect_0_program_memory_s1_clken)                           //                                         .clken
	);

	medidor_desempenho_irq_mapper irq_mapper (
		.clk           (clk_clk),                            //       clk.clk
		.reset         (rst_controller_001_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),           // receiver0.irq
		.sender_irq    (nios2_qsys_0_irq_irq)                //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                 // reset_in0.reset
		.clk            (clk_clk),                        //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.reset_in1      (nios2_qsys_0_debug_reset_request_reset), // reset_in1.reset
		.clk            (clk_clk),                                //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_001_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

endmodule
